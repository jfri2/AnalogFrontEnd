-------------------------------------------------------------------------------
-- <copyright_statement>
-- COPYRIGHT 2017 JOHN FRITZ. ALL RIGHTS RESERVED.
-- </copyright_statement>
--
-- <rights>
-- </rights>
--
-- <authors>
-- John Fritz
-- </authors>
--
-- <title>
-- interpolator.vhd
-- </title>
--
-- <description>
-- </description>
-------------------------------------------------------------------------------

--LIBRARY ieee;
--USE ieee.std_logic_1164.all;
--use ieee.numeric_std.all;
--
--ENTITY interpolator IS
--    PORT (
--
--    );
--END interpolator;
--
--ARCHITECTURE behavior OF interpolator IS
--
--BEGIN
--
--END behavior;
